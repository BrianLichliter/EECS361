-- This package is used for EECS 361 from Northwestern University.
-- by Kaicheng Zhang (kaichengz@gmail.com)

library ieee;
use ieee.std_logic_1164.all;
use work.eecs361_gates.all;

package eecs361 is
  -- Decoders
  component dec_n
    generic (
      -- Widths of the inputs.
      n	  : integer
    );
    port (
      src   : in std_logic_vector(n-1 downto 0);
      z	    : out std_logic_vector((2**n)-1 downto 0)
    );
  end component dec_n;

  -- Multiplexors
  component mux
    port (
      sel   : in  std_logic;
      src0  : in  std_logic;
      src1  : in  std_logic;
      z     : out std_logic
    );
  end component mux;

  component mux_n
    generic (
      -- Widths of the inputs.
      n	  : integer
    );
    port (
      sel   : in  std_logic;
      src0  : in  std_logic_vector(n-1 downto 0);
      src1  : in  std_logic_vector(n-1 downto 0);
      z     : out std_logic_vector(n-1 downto 0)
    );
  end component mux_n;

  component mux_32
    port (
      sel   : in  std_logic;
      src0  : in  std_logic_vector(31 downto 0);
      src1  : in  std_logic_vector(31 downto 0);
      z	    : out std_logic_vector(31 downto 0)
    );
  end component mux_32;

  component mux_1_4
    port (
      sel	: in  std_logic_vector(1 downto 0);
      src0	: in  std_logic;
      src1	: in  std_logic;
      src2	: in  std_logic;
      src3	: in  std_logic;
      z		: out std_logic
    );
  end component mux_1_4;

  component mux_n_4 is
    generic (
      n	: integer
    );
    port (
      sel  : in  std_logic_vector(1 downto 0);
      src0 : in  std_logic_vector(n-1 downto 0);
      src1 : in  std_logic_vector(n-1 downto 0);
      src2 : in  std_logic_vector(n-1 downto 0);
      src3 : in  std_logic_vector(n-1 downto 0);
      z    : out std_logic_vector(n-1 downto 0)
    );
  end component mux_n_4;

  -- Flip-flops

  -- D Flip-flops from Figure C.8.4 with a falling edge trigger.
  component dff
    port (
      clk   : in  std_logic;
      d	    : in  std_logic;
      q	    : out std_logic
    );
  end component dff;

  -- D Flip-flops from Figure C.8.4 with a rising edge trigger.
  component dffr
    port (
      clk   : in  std_logic;
      d	    : in  std_logic;
      q	    : out std_logic
    );
  end component dffr;

  -- D Flip-flops from Example 13-40 in http://www.altera.com/literature/hb/qts/qts_qii51007.pdf
  component dffr_a
    port (
      clk	 : in  std_logic;
      arst   : in  std_logic;
      aload  : in  std_logic;
      adata  : in  std_logic;
      d	     : in  std_logic;
      enable : in  std_logic;
      q	     : out std_logic
    );

  end component dffr_a;

  -- A 32bit SRAM from Figure C.9.1. It can only be used for simulation.
  component sram
	generic (
	  mem_file	: string
	);
	port (
	  -- chip select
	  cs	: in  std_logic;
	  -- output enable
	  oe	: in  std_logic;
	  -- write enable
	  we	: in  std_logic;
	  -- address line
	  addr	: in  std_logic_vector(31 downto 0);
	  -- data input
	  din	: in  std_logic_vector(31 downto 0);
	  -- data output
	  dout	: out std_logic_vector(31 downto 0)
	);
  end component sram;

  -- Synchronous SRAM with asynchronous reset.
  component syncram
    generic (
	  mem_file	: string
	);
	port (
      -- clock
      clk   : in  std_logic;
	  -- chip select
	  cs	: in  std_logic;
      -- output enable
	  oe	: in  std_logic;
	  -- write enable
	  we	: in  std_logic;
	  -- address line
	  addr	: in  std_logic_vector(31 downto 0);
	  -- data input
	  din	: in  std_logic_vector(31 downto 0);
	  -- data output
	  dout	: out std_logic_vector(31 downto 0)
	);
  end component syncram;

  -- n-bit full adder.
  component fulladder_n
    generic (
      n : integer
    );
    port (
      cin   : in std_logic;
      x     : in std_logic_vector(n-1 downto 0);
      y     : in std_logic_vector(n-1 downto 0);
      cout  : out std_logic;
      z     : out std_logic_vector(n-1 downto 0)
    );
  end component fulladder_n;

  -- 32-bit full adder.
  component fulladder_32
    port (
      cin   : in std_logic;
      x     : in std_logic_vector(31 downto 0);
      y     : in std_logic_vector(31 downto 0);
      z     : out std_logic_vector(31 downto 0);
      cout  : out std_logic
    );
  end component fulladder_32;

  -- 1-bit full adder.
  component fulladder_1
    port (
      x    : in std_logic;
      y    : in std_logic;
      cin  : in std_logic;
      z    : out std_logic;
      cout : out std_logic
    );
  end component fulladder_1;

  -- n-bit full adder.
  component fulladder_s_n
    generic (
      n : integer
    );
    port (
      A    : in std_logic_vector(n-1 downto 0);
      B    : in std_logic_vector(n-1 downto 0);
      R    : out std_logic_vector(n-1 downto 0)
    );
  end component fulladder_s_n;

  -- Cache tester.
  component cache_test
    generic (
      addr_trace_file : string;
      data_trace_file : string
    );
    port (
      DataIn : in std_logic_vector(31 downto 0);
      clk : in std_logic;
      Ready : in std_logic;
      rst : in std_logic;
      Addr : out std_logic_vector(31 downto 0);
      Data : out Std_logic_vector(31 downto 0);
      WR : out std_logic;
      Err : out std_logic
    );
  end component cache_test;

  -- Custom RAM
  component csram
    generic (
      INDEX_WIDTH : integer;
      BIT_WIDTH : integer
    );
    port (
      cs	  : in	std_logic;
      oe	  :	in	std_logic;
      we	  :	in	std_logic;
      index   : in	std_logic_vector(INDEX_WIDTH-1 downto 0);
      din	  :	in	std_logic_vector(BIT_WIDTH-1 downto 0);
      dout    :	out std_logic_vector(BIT_WIDTH-1 downto 0)
    );
  end component csram;

  component cmp_n
    generic (
      n : integer
    );
    port (
      a      : in std_logic_vector(n-1 downto 0);
      b      : in std_logic_vector(n-1 downto 0);

      a_eq_b : out std_logic;
      a_gt_b : out std_logic;
      a_lt_b : out std_logic;

      signed_a_gt_b : out std_logic;
      signed_a_lt_b : out std_logic
    );
  end component cmp_n;

  component comparator_1 is
    port (
      x   : in std_logic;
      y   : in std_logic;
      cin : in std_logic;
      z   : out std_logic
    );
  end component comparator_1;

  component comparator_32 is
    port (
      A   : in std_logic_vector(31 downto 0);
      B   : in std_logic_vector(31 downto 0);
      sgn : in std_logic; --1: signed compare, 0: unsigned compare
      R   : out std_logic_vector(31 downto 0) -- result
    );
  end component comparator_32;

  component ALU_1 is
    port (
      A    : in std_logic;
      B    : in std_logic;
      sel  : in std_logic_vector(1 downto 0);
      cin  : in std_logic;
      cout : out std_logic;
      R    : out std_logic
    );
  end component ALU_1;

  component ALU_32 is
    port (
      sel  : in std_logic_vector(1 downto 0);
      A    : in std_logic_vector(31 downto 0);
      B    : in std_logic_vector(31 downto 0);
      cin  : in std_logic;
      cout : out std_logic;  -- ?1? -> carry out
      ovf  : out std_logic;  -- ?1? -> overflow
      R    : out std_logic_vector(31 downto 0) -- result
    );
  end component ALU_32;

  component shifter_32 is
    port (
      A : in std_logic_vector(31 downto 0);
      B : in std_logic_vector(31 downto 0);
      R : out std_logic_vector(31 downto 0)
    );
  end component shifter_32;

  component signextender_n_m
    generic (
      n : integer;
      m : integer
    );
    port (
      A    : in std_logic_vector(n-1 downto 0);
      R    : out std_logic_vector(m-1 downto 0)
    );
  end component signextender_n_m;
  component and_5to1
      port (
          andIn : in std_logic_vector (4 downto 0);
          andOut : out std_logic
      );
  end component and_5to1;
  component decoder_5_32
     port (
         x : in std_logic_vector (4 downto 0);
         z : in std_logic_vector (31 downto 0)
     );
  end component decoder_5_32;
  component register_32bit
     port (
         clk : in std_logic;
       reset_active_low : in std_logic;
         write_en: in std_logic;
         D   : in std_logic_vector(31 downto 0);
         Z   : out std_logic_vector(31 downto 0)
     );
  end component register_32bit;

  component cpu
    generic (
      mem : string
    );
    port (
      clock   : in std_logic;
      reset   : in std_logic
    );
  end component cpu;

 component register_file
    port (
      clk : in std_logic;
      reset_active_low : in std_logic;
      write_en : in std_logic;
      write_data : in std_logic_vector(31 downto 0);
      read_index_A : in std_logic_vector(4 downto 0);
      read_index_B : in std_logic_vector(4 downto 0);
      write_index : in std_logic_vector(4 downto 0);
      read_op_A : out std_logic_vector(31 downto 0);
      read_op_B: out std_logic_vector(31 downto 0)
    );
 end component register_file;
 
 component control is 
     port ( 
  	   -- inputs from instruction
         opcode    : in  std_logic_vector(5 downto 0);
         func      : in  std_logic_vector(5 downto 0);
	     
	   -- 4 bit ALU control
         ALUCtr    : out std_logic_vector(3 downto 0);
   
	   -- 7 control signals
         regDst    : out std_logic;
         ALUSrc    : out std_logic;
         memtoReg  : out std_logic;
         regWrite  : out std_logic;
         memWrite  : out std_logic;
	       memRead	  : out std_logic;
         branch_eq    : out std_logic;
         branch_ne : out std_logic
     );
 end component control;
 
 component IFU is
   generic (
	   mem	: string
   );
   port (
	   clock	: in std_logic;
	   reset	: in std_logic;
	   branch_eq	: in std_logic;
	   branch_neq : in std_logic;
	   zero	: in std_logic;
	   inst	: inout std_logic_vector(31 downto 0)
   );
 end component IFU;
 
 component alu is
   port (
	   ctrl   : in std_logic_vector(3 downto 0);
	   A      : in std_logic_vector(31 downto 0);
	   B      : in std_logic_vector(31 downto 0);
	   cout   : out std_logic;  -- ?1? -> carry out
	   ovf    : out std_logic;  -- ?1? -> overflow
	   ze     : out std_logic;  -- ?1? -> is zero
	   R      : out std_logic_vector(31 downto 0) -- result
   );
 end component alu;
end;
